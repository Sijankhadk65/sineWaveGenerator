library ieee ;
use ieee.std_logic_1164.all;

entity CLK_E is
	port( 
		clk_o : OUT std_logic
	);
end entity CLK_E;

